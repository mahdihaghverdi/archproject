library ieee;
use ieee.std_logic_1164.all;

--  A testbench has no ports.
entity full_adder_tb is
end full_adder_tb;

architecture behav of full_adder_tb is
    --  Declaration of the component that will be instantiated.
    function to_string ( a: std_logic_vector) return string is
    variable b : string (1 to a'length) := (others => NUL);
    variable stri : integer := 1;
    begin
        for i in a'range loop
            b(stri) := std_logic'image(a((i)))(2);
        stri := stri+1;
        end loop;
    return b;
    end function;

    component full_adder
        port (
            a, b, ci : in std_logic_vector (31 downto 0);
            s, c : out std_logic_vector (31 downto 0)
        );
    end component;

    --  Specifies which entity is bound with the component.
    for full_adder_0: full_adder use entity work.full_adder;
    signal a, b, ci, s, c : std_logic_vector (31 downto 0);

begin
    --  Component instantiation.
    full_adder_0: full_adder port map (a => a, b => b, ci => ci, s => s, c => c);

--  This process does the real job.
process
    type pattern_type is record
        --  The inputs of the full_adder.
        a, b, ci : std_logic_vector (31 downto 0);
        --  The expected outputs of the full_adder.
        s, c : std_logic_vector (31 downto 0);
    end record;

--  The patterns to apply.
    type pattern_array is array (natural range <>) of pattern_type;
    constant patterns : pattern_array :=
        (
            (
                "00000100001110011000100011110101",
                "00000100001110011000100110100110",
                "00000000000000000000000000000000",
                "00000000000000000000000101010011",
                "00000100001110011000100010100100"
            ),
            (
                "01000100001110011010100011110101",
                "00111100001010111000000010100110",
                "00110111101111000010101001010010",
                "01001111101011100000001000000001",
                "00110100001110011010100011110110"
            ),
            (
                "11011100110111111011011011110100",
                "11100110111001101110101011011101",
                "10011110001001001010010111101110",
                "10100100000111011111100111000111",
                "11011110111001101010011011111100"
            ),
            (
                "01101000011010011100000011001000",
                "10010101010110100000010010000111",
                "11100011010000100000110000001101",
                "00011110011100011100100001000010",
                "11100001010010100000010010001101"
            ),
            (
                "00011010001011001100010110100111",
                "11101001011100010110010000101110",
                "01000100011101100111101011010110",
                "10110111001010111101101101011111",
                "01001000011101000110010010100110"
            ),
            (
                "11001010001100111000011100000010",
                "11110000101111010011111010011010",
                "11000101000011010010000000001000",
                "11111111100000111001100110010000",
                "11000000001111010010011000001010"
            ),
            (
                "00100110100011100101100100000111",
                "10101010110110011000011111001110",
                "01000010010101111111111111001101",
                "11001110000000000010000100000100",
                "00100010110111111101111111001111"
            ),
            (
                "11011101101111101100010110101111",
                "01001001111011001110110011010001",
                "10000100010011100101100111100110",
                "00010000000111000111000010011000",
                "11001101111011101100110111100111"
            ),
            (
                "11110001001000010001101001111100",
                "10001101000010100010100101100101",
                "10110111100010100001110111000110",
                "11001011101000010010111011011111",
                "10110101000010100001100101100100"
            ),
            (
                "11101011111010000110010010101011",
                "10101110010010000101110110011111",
                "00100110010111011110011100000010",
                "01100011111111011101111000110110",
                "10101110010010000110010110001011"
            ),
            (
                "01010010110000001100001111010111",
                "10010011100101111010001001110000",
                "00111011100111010001000010000111",
                "11111010110010100111000100100000",
                "00010011100101011000001011010111"
            ),
            (
                "10100100000111100110111100100100",
                "11101000100010100001101100111101",
                "01000100100111001011111100000011",
                "00001000000010001100101100011010",
                "11100100100111100011111100100101"
            ),
            (
                "10111111011011011001110001011011",
                "01000010111000000100111001010000",
                "11001000011000001100111000100011",
                "00110101111011010001110000101000",
                "11001010011000001100111001010011"
            ),
            (
                "01010000011011010100100110000100",
                "01110101110010001101100010000001",
                "11000111111111100111011111011001",
                "11100010010110111110011011011100",
                "01010101111011000101100110000001"
            ),
            (
                "00011010000101011110110110110100",
                "00000011000001100101010110010001",
                "00000011000011111001011100001101",
                "00011010000111000010111100101000",
                "00000011000001111101010110010101"
            ),
            (
                "01110101110101101101100011101001",
                "11001001001110110111111001101111",
                "00111000011100110100001001001101",
                "10000100100111101110010011001011",
                "01111001011100110101101001101101"
            ),
            (
                "01110001000101000101011000101001",
                "10101101000100010101111110100011",
                "01001111011001110000000011111100",
                "10010011011000100000100101110110",
                "01101101000101010101011010101001"
            ),
            (
                "01010101000001111011000110011100",
                "00010110110001000110010000001000",
                "01100101110101001000110010001000",
                "00100110000101110101100100011100",
                "01010101110001001010010010001000"
            ),
            (
                "10101100010010011001011101111011",
                "00101100111110100000000100001010",
                "00010000010100001000001000110100",
                "10010000111000110001010001000101",
                "00101100010110001000001100111010"
            ),
            (
                "01001010001111101011100001000010",
                "01100001001100100100100010111011",
                "10001011101100000001011111011001",
                "10100000101111001110011100100000",
                "01001011001100100001100011011011"
            ),
            (
                "10110101010100010110111010100010",
                "11100110101100111100110101001000",
                "10110111101110111101001110011111",
                "11100100010110010111000001110101",
                "10110111101100111100111110001010"
            ),
            (
                "01101001010101000100010110001100",
                "11010100010110110110100110111001",
                "10100101101010001011110000100000",
                "00011000101001111001000000010101",
                "11100101010110000110110110101000"
            ),
            (
                "11110101101111000110111010100101",
                "10111100010100100010111100101101",
                "11000011001001011101101111000100",
                "10001010110010111001101001001100",
                "11110101001101000110111110100101"
            ),
            (
                "01010101111110101010100011011100",
                "11110100111000010001010001100000",
                "01100111111111100111110010010010",
                "11000110111001011100000000101110",
                "01110101111110100011110011010000"
            )
        );

begin
    --  Check each pattern.
    for i in patterns'range loop
    --  Set the inputs.
    a <= patterns(i).a;
    b <= patterns(i).b;
    ci <= patterns(i).ci;
    --  Wait for the results.
    wait for 1 ns;
        --  Check the outputs.
            assert s = patterns(i).s
                report LF &
                "a : " & to_string(a) & LF &
                "b : " & to_string(b) & LF &
                "ci : " & to_string(ci) & LF &
                "s : " & to_string(s) & LF &
                "c : " & to_string(c) & LF &
                "Bad sum value";
            assert c = patterns(i).c
                report LF &
                "a : " & to_string(a) & LF &
                "b : " & to_string(b) & LF &
                "ci : " & to_string(ci) & LF &
                "s : " & to_string(s) & LF &
                "c : " & to_string(c) & LF &
                "Bad carry out value";
        end loop;
            assert false report "end of test" severity note;
        wait;
    end process;
end behav;
